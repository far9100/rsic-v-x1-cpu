// RISC-V 32IM CPU Testbench for Multiplication
// File: hardware/sim/tb_mul_test.v

`timescale 1ns / 1ps

module tb_mul_test;

    // Parameters
    localparam CLK_PERIOD = 10; // Clock period in ns (e.g., 100 MHz clock)
    localparam RESET_DURATION = CLK_PERIOD * 5; // How long to hold reset active
    localparam MAX_SIM_CYCLES = 500; // Maximum simulation cycles
    localparam MEM_SIZE_WORDS = 1024; // Memory size in words

    // Testbench signals
    reg         clk;
    reg         rst_n;

    // DUT (Device Under Test) Interface signals
    wire [31:0] i_mem_addr;
    reg  [31:0] i_mem_rdata; // Driven by testbench based on i_mem_addr

    wire [31:0] d_mem_addr;
    wire [31:0] d_mem_wdata;
    wire [3:0]  d_mem_wen;
    reg  [31:0] d_mem_rdata; // Driven by testbench based on d_mem_addr

    // Instantiate the CPU
    cpu_top u_cpu (
        .clk            (clk),
        .rst_n          (rst_n),
        .i_mem_addr     (i_mem_addr),
        .i_mem_rdata    (i_mem_rdata),
        .d_mem_addr     (d_mem_addr),
        .d_mem_wdata    (d_mem_wdata),
        .d_mem_wen      (d_mem_wen),
        .d_mem_rdata    (d_mem_rdata)
    );

    // Memory models (simplified)
    // Instruction Memory (ROM-like)
    reg [31:0] instr_mem [0:MEM_SIZE_WORDS-1];
    integer i;
    initial begin
        // Load instructions from a .hex file (e.g., generated by assembler)
        // IMPORTANT: Ensure this path is correct relative to where vvp is run (usually project root)
        $readmemh("tests/hex_outputs/mul_integrated_test.hex", instr_mem);
        
        // Initialize data memory (e.g., to zeros)
        for (i = 0; i < MEM_SIZE_WORDS; i = i + 1) begin
            data_mem[i] = 32'b0;
        end
    end

    // Instruction memory read logic (combinational)
    always @(*) begin
        if (i_mem_addr < 4*MEM_SIZE_WORDS) begin // Check bounds (byte address vs word array)
            i_mem_rdata = instr_mem[i_mem_addr / 4];
        end else begin
            i_mem_rdata = 32'hdeadbeef; // Out of bounds, return a recognizable invalid instruction
        end
    end

    // Data Memory (RAM-like)
    reg [31:0] data_mem [0:MEM_SIZE_WORDS-1];

    // Data memory read logic (combinational)
    always @(*) begin
        if (d_mem_addr < 4*MEM_SIZE_WORDS) begin // Check bounds
            d_mem_rdata = data_mem[d_mem_addr / 4];
        end else begin
            d_mem_rdata = 32'hxxxxxxxx; // Out of bounds
        end
    end

    // Data memory write logic (synchronous to clock)
    always @(posedge clk) begin
        if (rst_n) begin // Only write if not in reset
            if (d_mem_wen != 4'b0000 && d_mem_addr < 4*MEM_SIZE_WORDS) begin
                if (d_mem_wen == 4'b1111) begin // Word write
                    data_mem[d_mem_addr / 4] <= d_mem_wdata;
                    // Display memory writes for debugging
                    $display("DataMem Write: Addr=0x%h, Data=0x%h", d_mem_addr, d_mem_wdata);
                end
            end
        end
    end

    // Clock generation
    initial begin
        clk = 0;
        forever #(CLK_PERIOD / 2) clk = ~clk;
    end

    // Reset generation
    initial begin
        rst_n = 0; // Assert reset
        #(RESET_DURATION);
        rst_n = 1; // De-assert reset
    end

    // Simulation control and monitoring
    integer cycle_count_sim = 0;
    initial begin
        $display("Starting RISC-V CPU Multiplication Test Simulation...");
        wait (rst_n === 1);
        $display("Reset de-asserted. CPU operation begins at time %0t.", $time);

        for (cycle_count_sim = 0; cycle_count_sim < MAX_SIM_CYCLES; cycle_count_sim = cycle_count_sim + 1) begin
            @(posedge clk);
            // Print instruction being fetched every 50 cycles
            if (cycle_count_sim % 50 == 0) begin
                $display("Cycle %0d (sim): Fetching Instruction: %h", cycle_count_sim, i_mem_rdata);
            end
        end

        $display("Simulation finished at time %0t.", $time);
        $finish;
    end

    // Waveform dumping
    initial begin
        $dumpfile("tb_mul_test.vcd");
        $dumpvars(0, tb_mul_test);
    end

endmodule 