// RISC-V 32IM CPU Testbench
// File: hardware/sim/tb_cpu.v

`timescale 1ns / 1ps

module tb_cpu;

    // Parameters
    localparam CLK_PERIOD = 10; // Clock period in ns (e.g., 100 MHz clock)
    localparam RESET_DURATION = CLK_PERIOD * 5; // How long to hold reset active
    localparam MAX_SIM_CYCLES = 1000; // Maximum simulation cycles to prevent infinite run
    localparam MEM_SIZE_WORDS = 1024; // Memory size in words

    // Testbench signals
    reg         clk;
    reg         rst_n;

    // DUT (Device Under Test) Interface signals
    wire [31:0] i_mem_addr;
    reg  [31:0] i_mem_rdata; // Driven by testbench based on i_mem_addr

    wire [31:0] d_mem_addr;
    wire [31:0] d_mem_wdata;
    wire [3:0]  d_mem_wen;
    reg  [31:0] d_mem_rdata; // Driven by testbench based on d_mem_addr

    // Instantiate the CPU
    cpu_top u_cpu (
        .clk            (clk),
        .rst_n          (rst_n),
        .i_mem_addr     (i_mem_addr),
        .i_mem_rdata    (i_mem_rdata),
        .d_mem_addr     (d_mem_addr),
        .d_mem_wdata    (d_mem_wdata),
        .d_mem_wen      (d_mem_wen),
        .d_mem_rdata    (d_mem_rdata)
    );

    // Memory models (simplified)
    // Instruction Memory (ROM-like)
    reg [31:0] instr_mem [0:MEM_SIZE_WORDS-1];
    integer i;
    initial begin
        // Load instructions from a .hex file (e.g., generated by assembler)
        // IMPORTANT: Ensure this path is correct relative to where vvp is run (usually project root)
        $readmemh("tests/hex_outputs/add_test.hex", instr_mem);

        // The following hardcoded initialization is now REMOVED/COMMENTED
        // to ensure we use the .hex file.
        /*
        instr_mem[0] = 32'h00100113; // addi x2, x0, 1  (x2 = 1)
        instr_mem[1] = 32'h00200193; // addi x3, x0, 2  (x3 = 2)
        instr_mem[2] = 32'h00310233; // add  x4, x2, x3  (x4 = x2 + x3 = 3)
        instr_mem[3] = 32'h00000013; // NOP (addi x0, x0, 0) - to halt or observe
        
        // Ensure remaining memory is initialized, e.g. to NOP
        // This loop might not be necessary if $readmemh fills up to the program size
        // and the program ends with a halt, preventing execution of uninitialized memory.
        // However, for safety, or if $readmemh doesn't fill all, initialize to NOP.
        // This should ideally happen *after* $readmemh if $readmemh only partially fills.
        // For now, $readmemh is expected to handle the program part.
        // The warning "Not enough words" means $readmemh read fewer than MEM_SIZE_WORDS.
        // It's often better to initialize first, then $readmemh overwrites the start.
        for (i = 0; i < MEM_SIZE_WORDS; i = i + 1) begin
             instr_mem[i] = 32'h00000013; // Default to NOP
        end
        $readmemh("tests/hex_outputs/add_test.hex", instr_mem); // Read after default init
        */
    end

    // Instruction memory read logic (combinational)
    always @(*) begin
        if (i_mem_addr < 4*MEM_SIZE_WORDS) begin // Check bounds (byte address vs word array)
            i_mem_rdata = instr_mem[i_mem_addr / 4];
        end else begin
            i_mem_rdata = 32'hdeadbeef; // Out of bounds, return a recognizable invalid instruction
        end
    end

    // Data Memory (RAM-like)
    reg [31:0] data_mem [0:MEM_SIZE_WORDS-1];
    integer j;
    initial begin
        // Initialize data memory (e.g., to zeros)
        for (j = 0; j < MEM_SIZE_WORDS; j = j + 1) begin
            data_mem[j] = 32'b0;
        end
    end

    // Data memory read logic (combinational)
    always @(*) begin
        if (d_mem_addr < 4*MEM_SIZE_WORDS) begin // Check bounds
            d_mem_rdata = data_mem[d_mem_addr / 4];
        end else begin
            d_mem_rdata = 32'hxxxxxxxx; // Out of bounds
        end
    end

    // Data memory write logic (synchronous to clock)
    always @(posedge clk) begin
        if (rst_n) begin // Only write if not in reset
            if (d_mem_wen != 4'b0000 && d_mem_addr < 4*MEM_SIZE_WORDS) begin
                if (d_mem_wen == 4'b1111) begin // Word write
                    data_mem[d_mem_addr / 4] <= d_mem_wdata;
                    // Calculate cycle number relative to end of reset
                    // RESET_DURATION / CLK_PERIOD gives the number of reset cycles
                    // integer cycle_after_reset = ($time / CLK_PERIOD) - (RESET_DURATION / CLK_PERIOD);
                    // if (cycle_after_reset < 0) cycle_after_reset = 0; // Ensure non-negative during reset
                    // $display("Cycle %0d (eff): DataMem Write: Addr=0x%h, Data=0x%h", cycle_after_reset, d_mem_addr, d_mem_wdata);
                    $display("DataMem Write: Addr=0x%h, Data=0x%h", d_mem_addr, d_mem_wdata);
                end
            end
        end
    end

    // Clock generation
    initial begin
        clk = 0;
        forever #(CLK_PERIOD / 2) clk = ~clk;
    end

    // Reset generation
    initial begin
        rst_n = 0; // Assert reset
        #(RESET_DURATION);
        rst_n = 1; // De-assert reset
    end

    // Simulation control and monitoring
    integer cycle_count_sim = 0;
    initial begin
        $display("Starting RISC-V CPU Simulation...");
        wait (rst_n === 1);
        $display("Reset de-asserted. CPU operation begins at time %0t.", $time);

        for (cycle_count_sim = 0; cycle_count_sim < MAX_SIM_CYCLES; cycle_count_sim = cycle_count_sim + 1) begin
            @(posedge clk);
            // Check specific register value at a certain cycle count *after reset*
            // The $time might be large due to reset duration.
            // Let's use a counter that starts after reset.
            if (cycle_count_sim == 20) begin // Adjusted cycle count for NOPs, and to ensure WB of add x4
                 // Accessing hierarchical Verilog names can be simulator-dependent or tricky.
                 // A safer way is to output relevant signals from cpu_top or use $test$plusargs for checks.
                 // For now, assuming direct access works for iVerilog for debugging.
                 $display("Cycle %0d (sim): Reg x4 = %h (expected 3 for simple test with NOPs)", cycle_count_sim, u_cpu.u_id_stage.u_reg_file.registers[4]);
            end
        end

        if (cycle_count_sim == MAX_SIM_CYCLES) begin
            $display("Max simulation cycles reached (%0d).", MAX_SIM_CYCLES);
        end
        $display("Simulation finished at time %0t.", $time);
        $finish;
    end

    // Waveform dumping
    initial begin
        $dumpfile("tb_cpu.vcd");
        $dumpvars(0, tb_cpu);
    end

endmodule
