// RISC-V 32IM CPU Testbench
// File: hardware/sim/tb_cpu.v

`timescale 1ns / 1ps

module tb_cpu;

    // Parameters
    localparam CLK_PERIOD = 10; // Clock period in ns (e.g., 100 MHz clock)
    localparam RESET_DURATION = CLK_PERIOD * 5; // How long to hold reset active
    localparam MAX_SIM_CYCLES = 1000; // Maximum simulation cycles to prevent infinite run

    // Testbench signals
    reg         clk;
    reg         rst_n;

    // DUT (Device Under Test) Interface signals
    wire [31:0] i_mem_addr;
    reg  [31:0] i_mem_rdata; // Driven by testbench based on i_mem_addr

    wire [31:0] d_mem_addr;
    wire [31:0] d_mem_wdata;
    wire [3:0]  d_mem_wen;
    reg  [31:0] d_mem_rdata; // Driven by testbench based on d_mem_addr

    // Instantiate the CPU
    cpu_top u_cpu (
        .clk            (clk),
        .rst_n          (rst_n),
        .i_mem_addr     (i_mem_addr),
        .i_mem_rdata    (i_mem_rdata),
        .d_mem_addr     (d_mem_addr),
        .d_mem_wdata    (d_mem_wdata),
        .d_mem_wen      (d_mem_wen),
        .d_mem_rdata    (d_mem_rdata)
    );

    // Memory models (simplified)
    // Instruction Memory (ROM-like)
    reg [31:0] instr_mem [0:1023]; // Example: 1K words (4KB) instruction memory
    initial begin
        // Load instructions from a .hex file (e.g., generated by assembler)
        // $readmemh("path_to_your_instruction_hex_file.hex", instr_mem);
        // For now, fill with NOPs or a simple program
        instr_mem[0] = 32'h00100113; // addi x2, x0, 1  (x2 = 1)
        instr_mem[1] = 32'h00200193; // addi x3, x0, 2  (x3 = 2)
        instr_mem[2] = 32'h00310233; // add  x4, x2, x3  (x4 = x2 + x3 = 3)
        instr_mem[3] = 32'h00000013; // NOP (addi x0, x0, 0) - to halt or observe
        // ... fill more or use $readmemh
        // Ensure remaining memory is initialized, e.g. to NOP
        for (integer i = 4; i < 1024; i = i + 1) begin
            instr_mem[i] = 32'h00000013; // NOP
        end
    end

    // Instruction memory read logic (combinational)
    // Addresses are word addresses for this simple model (i_mem_addr is byte address)
    always @(*) begin
        if (i_mem_addr < 4*1024) begin // Check bounds
             // Divide by 4 for word addressing if i_mem_addr is byte address
            i_mem_rdata = instr_mem[i_mem_addr / 4];
        end else begin
            i_mem_rdata = 32'hxxxxxxxx; // Out of bounds
        end
    end

    // Data Memory (RAM-like)
    reg [31:0] data_mem [0:1023]; // Example: 1K words (4KB) data memory
    integer j;
    initial begin
        // Initialize data memory (e.g., to zeros)
        for (j = 0; j < 1024; j = j + 1) begin
            data_mem[j] = 32'b0;
        end
    end

    // Data memory read logic (combinational)
    always @(*) begin
        if (d_mem_addr < 4*1024) begin // Check bounds
            // Divide by 4 for word addressing if d_mem_addr is byte address
            d_mem_rdata = data_mem[d_mem_addr / 4];
        end else begin
            d_mem_rdata = 32'hxxxxxxxx; // Out of bounds
        end
    end

    // Data memory write logic (synchronous to clock)
    always @(posedge clk) begin
        if (rst_n) begin // Only write if not in reset
            if (d_mem_wen != 4'b0000 && d_mem_addr < 4*1024) begin // If write enabled and in bounds
                // Assuming word write for now (d_mem_wen == 4'b1111)
                // For byte/half-word writes, more complex logic is needed here based on d_mem_wen and d_mem_addr[1:0]
                if (d_mem_wen == 4'b1111) begin // Word write
                    data_mem[d_mem_addr / 4] <= d_mem_wdata;
                    $display("Cycle %0d: DataMem Write: Addr=0x%h, Data=0x%h", $time/CLK_PERIOD, d_mem_addr, d_mem_wdata);
                end
                // Add handling for byte/half-word writes if necessary
            end
        end
    end

    // Clock generation
    initial begin
        clk = 0;
        forever #(CLK_PERIOD / 2) clk = ~clk;
    end

    // Reset generation
    initial begin
        rst_n = 0; // Assert reset
        #(RESET_DURATION);
        rst_n = 1; // De-assert reset
    end

    // Simulation control and monitoring
    integer cycle_count = 0;
    initial begin
        $display("Starting RISC-V CPU Simulation...");
        // Wait for reset to de-assert
        wait (rst_n === 1);
        $display("Reset de-asserted. CPU operation begins.");

        // Monitor signals (example)
        // $monitor("Time: %0t, PC: %h, Instr: %h, d_mem_addr: %h, d_mem_wdata: %h, d_mem_wen: %b",
        //          $time, u_cpu.i_mem_addr, i_mem_rdata, d_mem_addr, d_mem_wdata, d_mem_wen);

        // Run for a certain number of cycles or until a specific condition
        for (cycle_count = 0; cycle_count < MAX_SIM_CYCLES; cycle_count = cycle_count + 1) begin
            @(posedge clk);
            // Check for a halt condition, e.g., specific instruction or PC value
            // if (u_cpu.i_mem_addr == 32'hSOME_HALT_ADDRESS) begin
            //     $display("Halt condition met at PC = %h. Simulation stopping.", u_cpu.i_mem_addr);
            //     break;
            // end
            if (cycle_count == 10) begin // Example: check a register after a few cycles
                 $display("Cycle %0d: Reg x4 = %h (expected 3 for simple test)", cycle_count, u_cpu.u_id_stage.u_reg_file.registers[4]);
            end
        end

        if (cycle_count == MAX_SIM_CYCLES) begin
            $display("Max simulation cycles reached (%0d).", MAX_SIM_CYCLES);
        end
        $display("Simulation finished at time %0t.", $time);
        $finish;
    end

    // Waveform dumping (optional, for tools like GTKWave)
    initial begin
        $dumpfile("tb_cpu.vcd");
        $dumpvars(0, tb_cpu); // Dump all signals in tb_cpu and below
    end

endmodule
